`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/09 10:03:44
// Design Name: 
// Module Name: RAM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//   Daddr，数据存储器地址输入端口
//   DataIn，数据存储器数据输入端口
//   DataOut，数据存储器数据输出端口
//   RD，数据存储器读控制信号，为0读
//   WR，数据存储器写控制信号，为0写



module Data_Memory_tb(
);

endmodule
